library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

library work;
use work.defines.all;

entity pac_textures is
	port(
		texture_id :  in integer range 0 to 9-1;
		x          :  in integer range 0 to 16-1;
		y          :  in integer range 0 to 16-1;
		ARGB       : out VGA_ARGB_t
	);
end pac_textures;

architecture RTL of pac_textures is 
	signal s_dataout : integer range 0 to 1;
	subtype t is integer range 0 to 1;
	type st is array (0 to (9*16*16)-1) of t;

	constant c_memory : st := ( 

															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,


															0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,

															-- text 2

															0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
															1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,

															-- text_3
															0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,

															--text 4

															0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,

															--text 5
															0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,
															
															--	text 6
															0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,

															--text 7

															0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,

															--text 8
															0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
															0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,
															0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,
															0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,
															0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,
															0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0);
begin

	s_dataout <= c_memory(((texture_id * 16 * 16) + x  + y*16));										  

	color_map : process(s_dataout)
	begin	
		if (s_dataout = 1) then
			ARGB <= "1" & "110";
		else
			ARGB <= "0" & "000";
		end if ;
	end process;

end;
